library IEEE;
use IEEE.STD_LOGIC_1164.all;
 -- type <new_type> is
--  record
--    <type_name>        : std_logic_vector( 7 downto 0);
--    <type_name>        : std_logic;
-- end record;
-- Declare constants
-- constant <constant_name>		: time := <time_unit> ns;
-- constant <constant_name>		: integer := <value;
-- Declare functions and procedure
-- function <function_name>  (signal <signal_name> : in <type_declaration>) return <type_declaration>;
-- procedure <procedure_name> (<type_declaration> <constant_name>	: in <type_declaration>);
package my_types_pkg is 
  constant n		: integer := 6;
  type array1 is array (0 to 323, 0 to 7) of integer;
  type array2 is array (0 to 7) of std_logic_vector(n-1 downto 0); 
  type array3 is array (0 to 647) of std_logic_vector(n-1 downto 0); 
  type array4 is array (0 to 6) of std_logic_vector(n-1 downto 0);
  type array5 is array (0 to 323) of std_logic;
constant row_weight :array5 := ('0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'1',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0',
																			'0');
constant col_position : array1 := (( 1 ,     109   ,  136  , 217   ,  298  , 326   ,  352 , 0 )
,( 2     , 110   , 137   , 218   , 299   , 327   , 353   , 0 )
,( 3     , 111   , 138   , 219   , 300   , 328   , 354   , 0 )
,( 4     , 112   , 139   , 220   , 301   , 329   , 355   , 0 )
,( 5     , 113   , 140   , 221   , 302   , 330   , 356   , 0 )
,( 6     , 114   , 141   , 222   , 303   , 331   , 357   , 0 )
,( 7     , 115   , 142   , 223   , 304   , 332   , 358   , 0 )
,( 8     , 116   , 143   , 224   , 305   , 333   , 359   , 0 )
,( 9     , 117   , 144   , 225   , 306   , 334   , 360   , 0 )
,( 10    , 118   , 145   , 226   , 307   , 335   , 361   , 0 )
,( 11    , 119   , 146   , 227   , 308   , 336   , 362   , 0 )
,( 12    , 120   , 147   , 228   , 309   , 337   , 363   , 0 )
,( 13    , 121   , 148   , 229   , 310   , 338   , 364   , 0 )
,( 14    , 122   , 149   , 230   , 311   , 339   , 365   , 0 )
,( 15    , 123   , 150   , 231   , 312   , 340   , 366   , 0 )
,( 16    , 124   , 151   , 232   , 313   , 341   , 367   , 0 )
,( 17    , 125   , 152   , 233   , 314   , 342   , 368   , 0 )
,( 18    , 126   , 153   , 234   , 315   , 343   , 369   , 0 )
,( 19    , 127   , 154   , 235   , 316   , 344   , 370   , 0 )
,( 20    , 128   , 155   , 236   , 317   , 345   , 371   , 0 )
,( 21    , 129   , 156   , 237   , 318   , 346   , 372   , 0 )
,( 22    , 130   , 157   , 238   , 319   , 347   , 373   , 0 )
,( 23    , 131   , 158   , 239   , 320   , 348   , 374   , 0 )
,( 24    , 132   , 159   , 240   , 321   , 349   , 375   , 0 )
,( 25    , 133   , 160   , 241   , 322   , 350   , 376   , 0 )
,( 26    , 134   , 161   , 242   , 323   , 351   , 377   , 0 )
,( 27    , 135   , 162   , 243   , 324   , 325   , 378   , 0 )
,( 23    , 28    , 126   , 163   , 190   , 229   , 352   , 379   )
,( 24    , 29    , 127   , 164   , 191   , 230   , 353   , 380   )
,( 25    , 30    , 128   , 165   , 192   , 231   , 354   , 381   )
,( 26    , 31    , 129   , 166   , 193   , 232   , 355   , 382   )
,( 27    , 32    , 130   , 167   , 194   , 233   , 356   , 383   )
,( 1     , 33    , 131   , 168   , 195   , 234   , 357   , 384   )
,( 2     , 34    , 132   , 169   , 196   , 235   , 358   , 385   )
,( 3     , 35    , 133   , 170   , 197   , 236   , 359   , 386   )
,( 4     , 36    , 134   , 171   , 198   , 237   , 360   , 387   )
,( 5     , 37    , 135   , 172   , 199   , 238   , 361   , 388   )
,( 6     , 38    , 109   , 173   , 200   , 239   , 362   , 389   )
,( 7     , 39    , 110   , 174   , 201   , 240   , 363   , 390   )
,( 8     , 40    , 111   , 175   , 202   , 241   , 364   , 391   )
,( 9     , 41    , 112   , 176   , 203   , 242   , 365   , 392   )
,( 10    , 42    , 113   , 177   , 204   , 243   , 366   , 393   )
,( 11    , 43    , 114   , 178   , 205   , 217   , 367   , 394   )
,( 12    , 44    , 115   , 179   , 206   , 218   , 368   , 395   )
,( 13    , 45    , 116   , 180   , 207   , 219   , 369   , 396   )
,( 14    , 46    , 117   , 181   , 208   , 220   , 370   , 397   )
,( 15    , 47    , 118   , 182   , 209   , 221   , 371   , 398   )
,( 16    , 48    , 119   , 183   , 210   , 222   , 372   , 399   )
,( 17    , 49    , 120   , 184   , 211   , 223   , 373   , 400   )
,( 18    , 50    , 121   , 185   , 212   , 224   , 374   , 401   )
,( 19    , 51    , 122   , 186   , 213   , 225   , 375   , 402   )
,( 20    , 52    , 123   , 187   , 214   , 226   , 376   , 403   )
,( 21    , 53    , 124   , 188   , 215   , 227   , 377   , 404   )
,( 22    , 54    , 125   , 189   , 216   , 228   , 378   , 405   )
,( 7     , 55    , 119   , 241   , 271   , 379   , 406   , 0 )
,( 8     , 56    , 120   , 242   , 272   , 380   , 407   , 0 )
,( 9     , 57    , 121   , 243   , 273   , 381   , 408   , 0 )
,( 10    , 58    , 122   , 217   , 274   , 382   , 409   , 0 )
,( 11    , 59    , 123   , 218   , 275   , 383   , 410   , 0 )
,( 12    , 60    , 124   , 219   , 276   , 384   , 411   , 0 )
,( 13    , 61    , 125   , 220   , 277   , 385   , 412   , 0 )
,( 14    , 62    , 126   , 221   , 278   , 386   , 413   , 0 )
,( 15    , 63    , 127   , 222   , 279   , 387   , 414   , 0 )
,( 16    , 64    , 128   , 223   , 280   , 388   , 415   , 0 )
,( 17    , 65    , 129   , 224   , 281   , 389   , 416   , 0 )
,( 18    , 66    , 130   , 225   , 282   , 390   , 417   , 0 )
,( 19    , 67    , 131   , 226   , 283   , 391   , 418   , 0 )
,( 20    , 68    , 132   , 227   , 284   , 392   , 419   , 0 )
,( 21    , 69    , 133   , 228   , 285   , 393   , 420   , 0 )
,( 22    , 70    , 134   , 229   , 286   , 394   , 421   , 0 )
,( 23    , 71    , 135   , 230   , 287   , 395   , 422   , 0 )
,( 24    , 72    , 109   , 231   , 288   , 396   , 423   , 0 )
,( 25    , 73    , 110   , 232   , 289   , 397   , 424   , 0 )
,( 26    , 74    , 111   , 233   , 290   , 398   , 425   , 0 )
,( 27 	 , 75	 , 112	 , 234	  , 291	 , 399	 , 426	 , 0 )
,( 1	 , 76	 , 113	 , 235	 , 292	 , 400	 , 427	 , 0 )
,( 2	 , 77	 , 114	 , 236	 , 293	 , 401	 , 428	 , 0 )
,( 3	 , 78	 , 115	 , 237	 , 294	 , 402	 , 429	 , 0 )
,( 4	 , 79	 , 116	 , 238	 , 295	 , 403	 , 430	 , 0 )
,( 5	 , 80	 , 117	 , 239	 , 296	 , 404	 , 431	 , 0 )
,( 6	 , 81	 , 118	 , 240	 , 297	 , 405	 , 432	 , 0 )
,( 3	 , 82	 , 129	 , 242	 , 244	 , 406	 , 433	 , 0 )
,( 4	 , 83	 , 130	 , 243	 , 245	 , 407	 , 434	 , 0 )
,( 5	 , 84	 , 131	 , 217	 , 246	 , 408	 , 435	 , 0 )
,( 6	 , 85	 , 132	 , 218	 , 247	 , 409	 , 436	 , 0 )
,( 7	 , 86	 , 133	 , 219	 , 248	 , 410	 , 437	 , 0 )
,( 8	 , 87	 , 134	 , 220	 , 249	 , 411	 , 438	 , 0 )
,( 9	 , 88	 , 135	 , 221	 , 250	 , 412	 , 439	 , 0 )
,( 10	 , 89	 , 109	 , 222	 , 251	 , 413	 , 440	 , 0 )
,( 11	 , 90	 , 110	 , 223	 , 252	 , 414	 , 441	 , 0 )
,( 12	 , 91	 , 111	 , 224	 , 253	 , 415	 , 442	 , 0 )
,( 13	 , 92	 , 112	 , 225	 , 254	 , 416	 , 443	 , 0 )
,( 14	 , 93	 , 113	 , 226	 , 255	 , 417	 , 444	 , 0 )
,( 15	 , 94	 , 114	 , 227	 , 256	 , 418	 , 445	 , 0 )
,( 16	 , 95	 , 115	 , 228	 , 257	 , 419	 , 446	 , 0 )
,( 17	 , 96	 , 116	 , 229	 , 258	 , 420	 , 447	 , 0 )
,( 18	 , 97	 , 117	 , 230	 , 259	 , 421	 , 448	 , 0 )
,( 19	 , 98	 , 118	 , 231	 , 260	 , 422	 , 449	 , 0 )
,( 20	 , 99	 , 119	 , 232	 , 261	 , 423	 , 450	 , 0 )
,( 21	 , 100	 , 120	 , 233	 , 262	 , 424	 , 451	 , 0 )
,( 22	 , 101	 , 121	 , 234	 , 263	 , 425	 , 452	 , 0 )
,( 23	 , 102	 , 122	 , 235	 , 264	 , 426	 , 453	 , 0 )
,( 24	 , 103	 , 123	 , 236	 , 265	 , 427	 , 454	 , 0 )
,( 25	 , 104	 , 124	 , 237	 , 266	 , 428	 , 455	 , 0 )
,( 26	 , 105	 , 125	 , 238	 , 267	 , 429	 , 456	 , 0 )
,( 27	 , 106	 , 126	 , 239	 , 268	 , 430	 , 457	 , 0 )
,( 1	 , 107	 , 127	 , 240	 , 269	 , 431	 , 458	 , 0 )
,( 2	 , 108	 , 128	 , 241	 , 270	 , 432	 , 459	 , 0 )
,( 24	 , 112	 , 217	 , 280	 , 309	 , 433	 , 460	 , 0 )
,( 25	 , 113	 , 218	 , 281	 , 310	 , 434	 , 461	 , 0 )
,( 26	 , 114	 , 219	 , 282	 , 311	 , 435	 , 462	 , 0 )
,( 27	 , 115	 , 220	 , 283	 , 312	 , 436	 , 463	 , 0 )
,( 1	 , 116	 , 221	 , 284	 , 313	 , 437	 , 464	 , 0 )
,( 2	 , 117	 , 222	 , 285	 , 314	 , 438	 , 465	 , 0 )
,( 3	 , 118	 , 223	 , 286	 , 315	 , 439	 , 466	 , 0 )
,( 4	 , 119	 , 224	 , 287	 , 316	 , 440	 , 467	 , 0 )
,( 5	 , 120	 , 225	 , 288	 , 317	 , 441	 , 468	 , 0 )
,( 6	 , 121	 , 226	 , 289	 , 318	 , 442	 , 469	 , 0 )
,( 7	 , 122	 , 227	 , 290	 , 319	 , 443	 , 470	 , 0 )
,( 8	 , 123	 , 228	 , 291	 , 320	 , 444	 , 471	 , 0 )
,( 9	 , 124	 , 229	 , 292	 , 321	 , 445	 , 472	 , 0 )
,( 10	 , 125	 , 230	 , 293	 , 322	 , 446	 , 473	 , 0 )
,( 11	 , 126	 , 231	 , 294	 , 323	 , 447	 , 474	 , 0 )
,( 12	 , 127	 , 232	 , 295	 , 324	 , 448	 , 475	 , 0 )
,( 13	 , 128	 , 233	 , 296	 , 298	 , 449	 , 476	 , 0 )
,( 14	 , 129	 , 234	 , 297	 , 299	 , 450	 , 477	 , 0 )
,( 15	 , 130	 , 235	 , 271	 , 300	 , 451	 , 478	 , 0 )
,( 16	 , 131	 , 236	 , 272	 , 301	 , 452	 , 479	 , 0 )
,( 17	 , 132	 , 237	 , 273	 , 302	 , 453	 , 480	 , 0 )
,( 18	 , 133	 , 238	 , 274	 , 303	 , 454	 , 481	 , 0 )
,( 19	 , 134	 , 239	 , 275	 , 304	 , 455	 , 482	 , 0 )
,( 20	 , 135	 , 240	 , 276	 , 305	 , 456	 , 483	 , 0 )
,( 21	 , 109	 , 241	 , 277	 , 306	 , 457	 , 484	 , 0 )
,( 22	 , 110	 , 242	 , 278	 , 307	 , 458	 , 485	 , 0 )
,( 23	 , 111	 , 243	 , 279	 , 308	 , 459	 , 486	 , 0 )
,( 25	 , 78	 , 83	 , 126	 , 166	 , 227	 , 460	 , 487	 )
,( 26	 , 79	 , 84	 , 127	 , 167	 , 228	 , 461	 , 488	 )
,( 27	 , 80	 , 85	 , 128	 , 168	 , 229	 , 462	 , 489	 )
,( 1	 , 81	 , 86	 , 129	 , 169	 , 230	 , 463	 , 490	 )
,( 2	 , 55	 , 87	 , 130	 , 170	 , 231	 , 464	 , 491	 )
,( 3	 , 56	 , 88	 , 131	 , 171	 , 232	 , 465	 , 492	 )
,( 4	 , 57	 , 89	 , 132	 , 172	 , 233	 , 466	 , 493	 )
,( 5	 , 58	 , 90	 , 133	 , 173	 , 234	 , 467	 , 494	 )
,( 6	 , 59	 , 91	 , 134	 , 174	 , 235	 , 468	 , 495	 )
,( 7	 , 60	 , 92	 , 135	 , 175	 , 236	 , 469	 , 496	 )
,( 8	 , 61	 , 93	 , 109	 , 176	 , 237	 , 470	 , 497	 )
,( 9	 , 62	 , 94	 , 110	 , 177	 , 238	 , 471	 , 498	 )
,( 10	 , 63	 , 95	 , 111	 , 178	 , 239	 , 472	 , 499	 )
,( 11	 , 64	 , 96	 , 112	 , 179	 , 240	 , 473	 , 500	 )
,( 12	 , 65	 , 97	 , 113	 , 180	 , 241	 , 474	 , 501	 )
,( 13	 , 66	 , 98	 , 114	 , 181	 , 242	 , 475	 , 502	 )
,( 14	 , 67	 , 99	 , 115	 , 182	 , 243	 , 476	 , 503	 )
,( 15	 , 68	 , 100	 , 116	 , 183	 , 217	 , 477	 , 504	 )
,( 16	 , 69	 , 101	 , 117	 , 184	 , 218	 , 478	 , 505	 )
,( 17	 , 70	 , 102	 , 118	 , 185	 , 219	 , 479	 , 506	 )
,( 18	 , 71	 , 103	 , 119	 , 186	 , 220	 , 480	 , 507	 )
,( 19	 , 72	 , 104	 , 120	 , 187	 , 221	 , 481	 , 508	 )
,( 20	 , 73	 , 105	 , 121	 , 188	 , 222	 , 482	 , 509	 )
,( 21	 , 74	 , 106	 , 122	 , 189	 , 223	 , 483	 , 510	 )
,( 22	 , 75	 , 107	 , 123	 , 163	 , 224	 , 484	 , 511	 )
,( 23	 , 76	 , 108	 , 124	 , 164	 , 225	 , 485	 , 512	 )
,( 24	 , 77	 , 82	 , 125	 , 165	 , 226	 , 486	 , 513	 )
,( 26	 , 117	 , 224	 , 262	 , 325	 , 487	 , 514	 , 0 )
,( 27	 , 118	 , 225	 , 263	 , 326	 , 488	 , 515	 , 0 )
,( 1	 , 119	 , 226	 , 264	 , 327	 , 489	 , 516	 , 0 )
,( 2	 , 120	 , 227	 , 265	 , 328	 , 490	 , 517	 , 0 )
,( 3	 , 121	 , 228	 , 266	 , 329	 , 491	 , 518	 , 0 )
,( 4	 , 122	 , 229	 , 267	 , 330	 , 492	 , 519	 , 0 )
,( 5	 , 123	 , 230	 , 268	 , 331	 , 493	 , 520	 , 0 )
,( 6	 , 124	 , 231	 , 269	 , 332	 , 494	 , 521	 , 0 )
,( 7	 , 125	 , 232	 , 270	 , 333	 , 495	 , 522	 , 0 )
,( 8	 , 126	 , 233	 , 244	 , 334	 , 496	 , 523	 , 0 )
,( 9	 , 127	 , 234	 , 245	 , 335	 , 497	 , 524	 , 0 )
,( 10	 , 128	 , 235	 , 246	 , 336	 , 498	 , 525	 , 0 )
,( 11	 , 129	 , 236	 , 247	 , 337	 , 499	 , 526	 , 0 )
,( 12	 , 130	 , 237	 , 248	 , 338	 , 500	 , 527	 , 0 )
,( 13	 , 131	 , 238	 , 249	 , 339	 , 501	 , 528	 , 0 )
,( 14	 , 132	 , 239	 , 250	 , 340	 , 502	 , 529	 , 0 )
,( 15	 , 133	 , 240	 , 251	 , 341	 , 503	 , 530	 , 0 )
,( 16	 , 134	 , 241	 , 252	 , 342	 , 504	 , 531	 , 0 )
,( 17	 , 135	 , 242	 , 253	 , 343	 , 505	 , 532	 , 0 )
,( 18	 , 109	 , 243	 , 254	 , 344	 , 506	 , 533	 , 0 )
,( 19	 , 110	 , 217	 , 255	 , 345	 , 507	 , 534	 , 0 )
,( 20	 , 111	 , 218	 , 256	 , 346	 , 508	 , 535	 , 0 )
,( 21	 , 112	 , 219	 , 257	 , 347	 , 509	 , 536	 , 0 )
,( 22	 , 113	 , 220	 , 258	 , 348	 , 510	 , 537	 , 0 )
,( 23	 , 114	 , 221	 , 259	 , 349	 , 511	 , 538	 , 0 )
,( 24	 , 115	 , 222	 , 260	 , 350	 , 512	 , 539	 , 0 )
,( 25	 , 116	 , 223	 , 261	 , 351	 , 513	 , 540	 , 0 )
,( 14	 , 52	 , 109	 , 171	 , 223	 , 514	 , 541	 , 0 )
,( 15	 , 53	 , 110	 , 172	 , 224	 , 515	 , 542	 , 0 )
,( 16	 , 54	 , 111	 , 173	 , 225	 , 516	 , 543	 , 0 )
,( 17	 , 28	 , 112	 , 174	 , 226	 , 517	 , 544	 , 0 )
,( 18	 , 29	 , 113	 , 175	 , 227	 , 518	 , 545	 , 0 )
,( 19	 , 30	 , 114	 , 176	 , 228	 , 519	 , 546	 , 0 )
,( 20	 , 31	 , 115	 , 177	 , 229	 , 520	 , 547	 , 0 )
,( 21	 , 32	 , 116	 , 178	 , 230	 , 521	 , 548	 , 0 )
,( 22	 , 33	 , 117	 , 179	 , 231	 , 522	 , 549	 , 0 )
,( 23	 , 34	 , 118	 , 180	 , 232	 , 523	 , 550	 , 0 )
,( 24	 , 35	 , 119	 , 181	 , 233	 , 524	 , 551	 , 0 )
,( 25	 , 36	 , 120	 , 182	 , 234	 , 525	 , 552	 , 0 )
,( 26	 , 37	 , 121	 , 183	 , 235	 , 526	 , 553	 , 0 )
,( 27	 , 38	 , 122	 , 184	 , 236	 , 527	 , 554	 , 0 )
,( 1	 , 39	 , 123	 , 185	 , 237	 , 528	 , 555	 , 0 )
,( 2	 , 40	 , 124	 , 186	 , 238	 , 529	 , 556	 , 0 )
,( 3	 , 41	 , 125	 , 187	 , 239	 , 530	 , 557	 , 0 )
,( 4	 , 42	 , 126	 , 188	 , 240	 , 531	 , 558	 , 0 )
,( 5	 , 43	 , 127	 , 189	 , 241	 , 532	 , 559	 , 0 )
,( 6	 , 44	 , 128	 , 163	 , 242	 , 533	 , 560	 , 0 )
,( 7	 , 45	 , 129	 , 164	 , 243	 , 534	 , 561	 , 0 )
,( 8	 , 46	 , 130	 , 165	 , 217	 , 535	 , 562	 , 0 )
,( 9	 , 47	 , 131	 , 166	 , 218	 , 536	 , 563	 , 0 )
,( 10	 , 48	 , 132	 , 167	 , 219	 , 537	 , 564	 , 0 )
,( 11	 , 49	 , 133	 , 168	 , 220	 , 538	 , 565	 , 0 )
,( 12	 , 50	 , 134	 , 169	 , 221	 , 539	 , 566	 , 0 )
,( 13	 , 51	 , 135	 , 170	 , 222	 , 540	 , 567	 , 0 )
,( 8	 , 48	 , 98	 , 131	 , 146	 , 240	 , 541	 , 568	 )
,( 9	 , 49	 , 99	 , 132	 , 147	 , 241	 , 542	 , 569	 )
,( 10	 , 50	 , 100	 , 133	 , 148	 , 242	 , 543	 , 570	 )
,( 11	 , 51	 , 101	 , 134	 , 149	 , 243	 , 544	 , 571	 )
,( 12	 , 52	 , 102	 , 135	 , 150	 , 217	 , 545	 , 572	 )
,( 13	 , 53	 , 103	 , 109	 , 151	 , 218	 , 546	 , 573	 )
,( 14	 , 54	 , 104	 , 110	 , 152	 , 219	 , 547	 , 574	 )
,( 15	 , 28	 , 105	 , 111	 , 153	 , 220	 , 548	 , 575	 )
,( 16	 , 29	 , 106	 , 112	 , 154	 , 221	 , 549	 , 576	 )
,( 17	 , 30	 , 107	 , 113	 , 155	 , 222	 , 550	 , 577	 )
,( 18	 , 31	 , 108	 , 114	 , 156	 , 223	 , 551	 , 578	 )
,( 19	 , 32	 , 82	 , 115	 , 157	 , 224	 , 552	 , 579	 )
,( 20	 , 33	 , 83	 , 116	 , 158	 , 225	 , 553	 , 580	 )
,( 21	 , 34	 , 84	 , 117	 , 159	 , 226	 , 554	 , 581	 )
,( 22	 , 35	 , 85	 , 118	 , 160	 , 227	 , 555	 , 582	 )
,( 23	 , 36	 , 86	 , 119	 , 161	 , 228	 , 556	 , 583	 )
,( 24	 , 37	 , 87	 , 120	 , 162	 , 229	 , 557	 , 584	 )
,( 25	 , 38	 , 88	 , 121	 , 136	 , 230	 , 558	 , 585	 )
,( 26	 , 39	 , 89	 , 122	 , 137	 , 231	 , 559	 , 586	 )
,( 27	 , 40	 , 90	 , 123	 , 138	 , 232	 , 560	 , 587	 )
,( 1	 , 41	 , 91	 , 124	 , 139	 , 233	 , 561	 , 588	 )
,( 2	 , 42	 , 92	 , 125	 , 140	 , 234	 , 562	 , 589	 )
,( 3	 , 43	 , 93	 , 126	 , 141	 , 235	 , 563	 , 590	 )
,( 4	 , 44	 , 94	 , 127	 , 142	 , 236	 , 564	 , 591	 )
,( 5	 , 45	 , 95	 , 128	 , 143	 , 237	 , 565	 , 592	 )
,( 6	 , 46	 , 96	 , 129	 , 144	 , 238	 , 566	 , 593	 )
,( 7	 , 47	 , 97	 , 130	 , 145	 , 239	 , 567	 , 594	 )
,( 12	 , 128	 , 230	 , 274	 , 315	 , 568	 , 595	 , 0 )
,( 13	 , 129	 , 231	 , 275	 , 316	 , 569	 , 596	 , 0 )
,( 14	 , 130	 , 232	 , 276	 , 317	 , 570	 , 597	 , 0 )
,( 15	 , 131	 , 233	 , 277	 , 318	 , 571	 , 598	 , 0 )
,( 16	 , 132	 , 234	 , 278	 , 319	 , 572	 , 599	 , 0 )
,( 17	 , 133	 , 235	 , 279	 , 320	 , 573	 , 600	 , 0 )
,( 18	 , 134	 , 236	 , 280	 , 321	 , 574	 , 601	 , 0 )
,( 19	 , 135	 , 237	 , 281	 , 322	 , 575	 , 602	 , 0 )
,( 20	 , 109	 , 238	 , 282	 , 323	 , 576	 , 603	 , 0 )
,( 21	 , 110	 , 239	 , 283	 , 324	 , 577	 , 604	 , 0 )
,( 22	 , 111	 , 240	 , 284	 , 298	 , 578	 , 605	 , 0 )
,( 23	 , 112	 , 241	 , 285	 , 299	 , 579	 , 606	 , 0 )
,( 24	 , 113	 , 242	 , 286	 , 300	 , 580	 , 607	 , 0 )
,( 25	 , 114	 , 243	 , 287	 , 301	 , 581	 , 608	 , 0 )
,( 26	 , 115	 , 217	 , 288	 , 302	 , 582	 , 609	 , 0 )
,( 27	 , 116	 , 218	 , 289	 , 303	 , 583	 , 610	 , 0 )
,( 1	 , 117	 , 219	 , 290	 , 304	 , 584	 , 611	 , 0 )
,( 2	 , 118	 , 220	 , 291	 , 305	 , 585	 , 612	 , 0 )
,( 3	 , 119	 , 221	 , 292	 , 306	 , 586	 , 613	 , 0 )
,( 4	 , 120	 , 222	 , 293	 , 307	 , 587	 , 614	 , 0 )
,( 5	 , 121	 , 223	 , 294	 , 308	 , 588	 , 615	 , 0 )
,( 6	 , 122	 , 224	 , 295	 , 309	 , 589	 , 616	 , 0 )
,( 7	 , 123	 , 225	 , 296	 , 310	 , 590	 , 617	 , 0 )
,( 8	 , 124	 , 226	 , 297	 , 311	 , 591	 , 618	 , 0 )
,( 9	 , 125	 , 227	 , 271	 , 312	 , 592	 , 619	 , 0 )
,( 10	 , 126	 , 228	 , 272	 , 313	 , 593	 , 620	 , 0 )
,( 11	 , 127	 , 229	 , 273	 , 314	 , 594	 , 621	 , 0 )
,( 26	 , 63	 , 132	 , 154	 , 204	 , 226	 , 595	 , 622	 )
,( 27	 , 64	 , 133	 , 155	 , 205	 , 227	 , 596	 , 623	 )
,( 1	 , 65	 , 134	 , 156	 , 206	 , 228	 , 597	 , 624	 )
,( 2	 , 66	 , 135	 , 157	 , 207	 , 229	 , 598	 , 625	 )
,( 3	 , 67	 , 109	 , 158	 , 208	 , 230	 , 599	 , 626	 )
,( 4	 , 68	 , 110	 , 159	 , 209	 , 231	 , 600	 , 627	 )
,( 5	 , 69	 , 111	 , 160	 , 210	 , 232	 , 601	 , 628	 )
,( 6	 , 70	 , 112	 , 161	 , 211	 , 233	 , 602	 , 629	 )
,( 7	 , 71	 , 113	 , 162	 , 212	 , 234	 , 603	 , 630	 )
,( 8	 , 72	 , 114	 , 136	 , 213	 , 235	 , 604	 , 631	 )
,( 9	 , 73	 , 115	 , 137	 , 214	 , 236	 , 605	 , 632	 )
,( 10	 , 74	 , 116	 , 138	 , 215	 , 237	 , 606	 , 633	 )
,( 11	 , 75	 , 117	 , 139	 , 216	 , 238	 , 607	 , 634	 )
,( 12	 , 76	 , 118	 , 140	 , 190	 , 239	 , 608	 , 635	 )
,( 13	 , 77	 , 119	 , 141	 , 191	 , 240	 , 609	 , 636	 )
,( 14	 , 78	 , 120	 , 142	 , 192	 , 241	 , 610	 , 637	 )
,( 15	 , 79	 , 121	 , 143	 , 193	 , 242	 , 611	 , 638	 )
,( 16	 , 80	 , 122	 , 144	 , 194	 , 243	 , 612	 , 639	 )
,( 17	 , 81	 , 123	 , 145	 , 195	 , 217	 , 613	 , 640	 )
,( 18	 , 55	 , 124	 , 146	 , 196	 , 218	 , 614	 , 641	 )
,( 19	 , 56	 , 125	 , 147	 , 197	 , 219	 , 615	 , 642	 )
,( 20	 , 57	 , 126	 , 148	 , 198	 , 220	 , 616	 , 643	 )
,( 21	 , 58	 , 127	 , 149	 , 199	 , 221	 , 617	 , 644	 )
,( 22	 , 59	 , 128	 , 150	 , 200	 , 222	 , 618	 , 645	 )
,( 23	 , 60	 , 129	 , 151	 , 201	 , 223	 , 619	 , 646	 )
,( 24	 , 61	 , 130	 , 152	 , 202	 , 224	 , 620	 , 647	 )
,( 25	 , 62	 , 131	 , 153	 , 203	 , 225	 , 621	 , 648	 )
,( 4	 , 125	 , 192	 , 242	 , 249	 , 326	 , 622	 , 0 )
,( 5	 , 126	 , 193	 , 243	 , 250	 , 327	 , 623	 , 0 )
,( 6	 , 127	 , 194	 , 217	 , 251	 , 328	 , 624	 , 0 )
,( 7	 , 128	 , 195	 , 218	 , 252	 , 329	 , 625	 , 0 )
,( 8	 , 129	 , 196	 , 219	 , 253	 , 330	 , 626	 , 0 )
,( 9	 , 130	 , 197	 , 220	 , 254	 , 331	 , 627	 , 0 )
,( 10	 , 131	 , 198	 , 221	 , 255	 , 332	 , 628	 , 0 )
,( 11	 , 132	 , 199	 , 222	 , 256	 , 333	 , 629	 , 0 )
,( 12	 , 133	 , 200	 , 223	 , 257	 , 334	 , 630	 , 0 )
,( 13	 , 134	 , 201	 , 224	 , 258	 , 335	 , 631	 , 0 )
,( 14	 , 135	 , 202	 , 225	 , 259	 , 336	 , 632	 , 0 )
,( 15	 , 109	 , 203	 , 226	 , 260	 , 337	 , 633	 , 0 )
,( 16	 , 110	 , 204	 , 227	 , 261	 , 338	 , 634	 , 0 )
,( 17	 , 111	 , 205	 , 228	 , 262	 , 339	 , 635	 , 0 )
,( 18	 , 112	 , 206	 , 229	 , 263	 , 340	 , 636	 , 0 )
,( 19	 , 113	 , 207	 , 230	 , 264	 , 341	 , 637	 , 0 )
,( 20	 , 114	 , 208	 , 231	 , 265	 , 342	 , 638	 , 0 )
,( 21	 , 115	 , 209	 , 232	 , 266	 , 343	 , 639	 , 0 )
,( 22	 , 116	 , 210	 , 233	 , 267	 , 344	 , 640	 , 0 )
,( 23	 , 117	 , 211	 , 234	 , 268	 , 345	 , 641	 , 0 )
,( 24	 , 118	 , 212	 , 235	 , 269	 , 346	 , 642	 , 0 )
,( 25	 , 119	 , 213	 , 236	 , 270	 , 347	 , 643	 , 0 )
,( 26	 , 120	 , 214	 , 237	 , 244	 , 348	 , 644	 , 0 )
,( 27	 , 121	 , 215	 , 238	 , 245	 , 349	 , 645	 , 0 )
,( 1	 , 122	 , 216	 , 239	 , 246	 , 350	 , 646	 , 0 )
,( 2	 , 123	 , 190	 , 240	 , 247	 , 351	 , 647	 , 0 )
,( 3	 , 124	 , 191	 , 241	 , 248	 , 325	 , 648	 , 0 ));

end my_types_pkg;

package body my_types_pkg is

---- Example 1
--  function <function_name>  (signal <signal_name> : in <type_declaration>  ) return <type_declaration> is
--    variable <variable_name>     : <type_declaration>;
--  begin
--    <variable_name> := <signal_name> xor <signal_name>;
--    return <variable_name>; 
--  end <function_name>;

---- Example 2
--  function <function_name>  (signal <signal_name> : in <type_declaration>;
--                         signal <signal_name>   : in <type_declaration>  ) return <type_declaration> is
--  begin
--    if (<signal_name> = '1') then
--      return <signal_name>;
--    else
--      return 'Z';
--    end if;
--  end <function_name>;

---- Procedure Example
--  procedure <procedure_name>  (<type_declaration> <constant_name>  : in <type_declaration>) is
--    
--  begin
--    
--  end <procedure_name>;
 
end my_types_pkg;
